library verilog;
use verilog.vl_types.all;
entity problem4tb is
end problem4tb;
