library verilog;
use verilog.vl_types.all;
entity pipeline_cpu_tb is
end pipeline_cpu_tb;
