library verilog;
use verilog.vl_types.all;
entity reg_32_tb is
end reg_32_tb;
