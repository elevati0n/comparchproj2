library verilog;
use verilog.vl_types.all;
entity problem5tb is
end problem5tb;
