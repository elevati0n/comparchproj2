library verilog;
use verilog.vl_types.all;
entity problem6tb is
end problem6tb;
