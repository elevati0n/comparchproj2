library verilog;
use verilog.vl_types.all;
entity test_mux2_1 is
end test_mux2_1;
